`include "uart_rx_config.sv"
`include "seq_item.sv"
`include "base_seq.sv"
`include "uart_rx_sequencer.sv"
`include "uart_rx_drv.sv"
`include "uart_rx_moni_in.sv"
`include "uart_rx_moni_out.sv"
`include "uart_rx_agent.sv"
`include "uart_rx_sb.sv"
`include "uart_rx_env.sv"
	